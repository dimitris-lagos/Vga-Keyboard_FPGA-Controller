module top(reset,clk,ps2clk,ps2data,hsync,vsync, Red, Green, Blue);input reset,clk;input ps2clk,ps2data;output hsync,vsync;output [2:0]Red,Green,Blue;wire [7:0]scancode,data_out;wire clkdiv4,display_area,clk,reset,flag,char_enable;wire [5:0] start_address_out,address_output;wire one_bit_output,r,g,b,fv;wire [3:0]line;wire[2:0] r1,g1,b1,up;pix_clk pix (clk,reset,clkdiv4);kbd_protocol kbdp (reset, clkdiv4, ps2clk, ps2data, scancode,flag);kbd_decoder kbdd (clkdiv4,reset,flag,scancode,start_address_out,r,g,b,fv,up,char_enable); vgasync syn (clk,clkdiv4,reset,up,hsync,vsync,display_area,line);iterator ite(line,display_area,start_address_out,address_output);char_rom chr (char_enable,address_output,data_out);shifter shf (reset,data_out,clkdiv4,display_area,one_bit_output);coloriser clr (reset,clk,clkdiv4,display_area,one_bit_output,r,g,b,r1,g1,b1);bonus bns (clkdiv4,reset,fv,vsync,r1,g1,b1,Red,Green,Blue);        endmodule 